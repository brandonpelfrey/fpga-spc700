module DSPVoice (
  
);
  
endmodule